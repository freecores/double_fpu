
`timescale 1ps / 1ps
module fpu_tb;


//Internal signals declarations:
reg clk;
reg rst;
reg enable;
reg fpu_op;
reg [63:0]opa;
reg [63:0]opb;
wire [63:0]out;
wire ready; 


	fpu UUT (
		.clk(clk),
		.rst(rst),
		.enable(enable),
		.fpu_op(fpu_op),
		.opa(opa),
		.opb(opb),
		.out(out),
		.ready(ready));

initial
begin : STIMUL 
	#0 
	enable = 1'b0;
	rst = 1'b1;
	fpu_op = 1'b1;
    #10000; //0
	enable = 1'b1;
	rst = 1'b0;	 
//inputA:-8.7700000000e+000
//inputB:4.9600000000e+000
opa = 64'b1100000000100001100010100011110101110000101000111101011100001010;
opb = 64'b0100000000010011110101110000101000111101011100001010001111010111;
fpu_op = 1'b0;
#10000;

//inputA:5.6668000000e+004
//inputB:2.3300000000e+002
opa = 64'b0100000011101011101010111000000000000000000000000000000000000000;
opb = 64'b0100000001101101001000000000000000000000000000000000000000000000;	   
fpu_op = 1'b1;		   
#10000;
//inputA:4.8999000000e+004
//inputB:3.4700000000e+001		
opa = 64'b0100000011100111111011001110000000000000000000000000000000000000;
opb = 64'b0100000001000001010110011001100110011001100110011001100110011010;
fpu_op = 1'b0;
#10000;

//inputA:1.0000000000e-200
//inputB:4.0000000000e-198
opa = 64'b0001011001101000011111101001001000010101010011101111011110101100;
opb = 64'b0001011011110011001000101110001000100000101001011011000101111110;
fpu_op = 1'b1;

#10000;
//inputA:8.9990000000e+003
//inputB:2.0000000000e-002
opa = 64'b0100000011000001100100111000000000000000000000000000000000000000;
opb = 64'b0011111110010100011110101110000101000111101011100001010001111011;
fpu_op = 1'b1;

#10000;
//inputA:4.4500000000e+002
//inputB:4.4437000000e+002
opa = 64'b0100000001111011110100000000000000000000000000000000000000000000;
opb = 64'b0100000001111011110001011110101110000101000111101011100001010010;
fpu_op = 1'b1;

#10000;	
//inputA:4.9342000000e+001
//inputB:2.3000000000e-002
opa = 64'b0100000001001000101010111100011010100111111011111001110110110010;
opb = 64'b0011111110010111100011010100111111011111001110110110010001011010;
fpu_op = 1'b0;


#10000;
//inputA:6.9100000000e+001
//inputB:6.8770000000e+001
opa = 64'b0100000001010001010001100110011001100110011001100110011001100110;
opb = 64'b0100000001010001001100010100011110101110000101000111101011100001;
fpu_op = 1'b0;

#10000;
//inputA:-8.9990000000e+003
//inputB:-9.5666000000e+004
opa = 64'b1100000011000001100100111000000000000000000000000000000000000000;
opb = 64'b1100000011110111010110110010000000000000000000000000000000000000;
fpu_op = 1'b0;

#10000;
//inputA:9.8300000000e+001
//inputB:-9.5666700000e+004
opa = 64'b0100000001011000100100110011001100110011001100110011001100110011;
opb = 64'b1100000011110111010110110010101100110011001100110011001100110011;
fpu_op = 1'b1;

#10000;
//inputA:6.8700000000e+001
//inputB:-9.5511000000e+002
opa = 64'b0100000001010001001011001100110011001100110011001100110011001101;
opb = 64'b1100000010001101110110001110000101000111101011100001010001111011;
fpu_op = 1'b0;

#10000;	   
//inputA:-9.5400000000e+001
//inputB:9.8100000000e+001
opa = 64'b1100000001010111110110011001100110011001100110011001100110011010;
opb = 64'b0100000001011000100001100110011001100110011001100110011001100110;
fpu_op = 1'b1;

#10000;	 
//inputA:-9.6300000000e+001
//inputB:9.8300000000e+001
opa = 64'b1100000001011000000100110011001100110011001100110011001100110011;
opb = 64'b0100000001011000100100110011001100110011001100110011001100110011;
fpu_op = 1'b0;

#10000;	 
//inputA:-4.5600000000e+001
//inputB:-9.8660000000e+001
opa = 64'b1100000001000110110011001100110011001100110011001100110011001101;
opb = 64'b1100000001011000101010100011110101110000101000111101011100001010;
fpu_op = 1'b1;

#10000;	
//inputA:2.0000000000e-308
//inputB:4.0000000000e-300
opa = 64'b0000000000001110011000011010110011110000001100111101000110100100;
opb = 64'b0000000111000101011011100001111111000010111110001111001101011001;
fpu_op = 1'b0;

#10000;	
//inputA:1.#INF000000e+000
//inputB:3.0000000000e+100
opa = 64'b0111111111110000000000000000000000000000000000000000000000000000;
opb = 64'b0101010011001011011011101000001110111000010111110010010100111011;
fpu_op = 1'b1;

#30000;		 
//Output:-3.810000000000000e+000
if (out==64'hC00E7AE147AE147C)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! C00E7AE147AE147C out is %h", out);
//Output:5.643500000000000e+004	
#10000;
if (out==64'h40EB8E6000000000)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 40EB8E6000000000 out is %h", out); 	
#10000;
	//Output:4.903370000000000e+004
if (out==64'h40E7F13666666666)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 40E7F13666666666 out is %h", out); 
#10000;
//Output:-3.990000000000000e-198
if (out==64'h96F316A2D79B0A03)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 96F316A2D79B0A03 out is %h", out);
#10000;
//Output:8.998980000000000e+003
if (out==64'h40C1937D70A3D70B)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 40C1937D70A3D70B out is %h", out);

#10000;
//Output:6.299999999999955e-001
if (out==64'h3FE428F5C28F5C00)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 3FE428F5C28F5C00 out is %h", out);


#10000;
//Output:4.936500000000000e+001
if (out==64'h4048AEB851EB851E)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 4048AEB851EB851E out is %h", out);

#10000;
//Output:1.378700000000000e+002
if (out==64'h40613BD70A3D70A3)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 40613BD70A3D70A3 out is %h", out);


#10000;
//Output:-1.046650000000000e+005
if (out==64'hC0F98D9000000000)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! C0F98D9000000000 out is %h", out);

#10000;
//Output:9.576500000000000e+004
if (out==64'h40F7614FFFFFFFFF)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 40F7614FFFFFFFFF out is %h", out);
 

#10000;
//Output:-8.864100000000001e+002
if (out==64'hC08BB347AE147AE2)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! C08BB347AE147AE2 out is %h", out);

#10000;
//Output:-1.935000000000000e+002
if (out==64'hC068300000000000)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! C068300000000000 out is %h", out);
 

#10000;
//Output:2.000000000000000e+000
if (out==64'h4000000000000000)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 4000000000000000 out is %h", out);

#10000;
//Output:5.306000000000000e+001
if (out==64'h404A87AE147AE148)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 404A87AE147AE148 out is %h", out);
 

#10000;
//Output:4.000000000000000e-300
if (out==64'h01C56E1FC2F8F359)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 01C56E1FC2F8F359 out is %h", out);

#10000;
//Output:1.#INF00000000000e+000
if (out==64'h7FF0000000000000)
	$display($time,"ps Answer is correct %h", out);
else
	$display($time,"ps Error! 7FF0000000000000 out is %h", out);

	
	#290000; 
	$finish;	
end 
	
always
begin : CLOCK_clk
	clk = 1'b0;
	#5000; 
	clk = 1'b1;
	#5000; 
end


endmodule
